-- Intentionally redacted